
module tb;
    initial begin
        #1;
        $finish();
    end
endmodule
